module cla_8bits(a,b,c0,c8,s);
input     [7:0]       a,b;
input                 c0;
output                c8;
output    [7:0]       s;
reg       [7:0]       p,q;
reg       [7:1]       c;
reg       [7:0]       s;
reg                   c8;
always@(a or b or c0)
begin
         p=a|b;
         q=a&b;
         
         c[1]=q[0]  |  p[0]&c0;
         c[2]=q[1]  |  p[1]&q[0]  |  p[1]&p[0]&c0;
         c[3]=q[2]  |  p[2]&q[1]  |  p[2]&p[1]&q[0]  |  p[2]&p[1]&p[0]&c0;
         c[4]=q[3]  |  p[3]&q[2]  |  p[3]&p[2]&q[1]  |  p[3]&p[2]&p[1]&q[0]  |  p[3]&p[2]&p[1]&p[0]&c0;
         c[5]=q[4]  |  p[4]&q[3]  |  p[4]&p[3]&q[2]  |  p[4]&p[3]&p[2]&q[1]  |  p[4]&p[3]&p[2]&p[1]&q[0]  |  p[4]&p[3]&p[2]&p[1]&p[0]&c0;
         c[6]=q[5]  |  p[5]&q[4]  |  p[5]&p[4]&q[3]  |  p[5]&p[4]&p[3]&q[2]  |  p[5]&p[4]&p[3]&p[2]&q[1]  |  p[5]&p[4]&p[3]&p[2]&p[1]&q[0]  |  p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c0;
         c[7]=q[6]  |  p[6]&q[5]  |  p[6]&p[5]&q[4]  |  p[6]&p[5]&p[4]&q[3]  |  p[6]&p[5]&p[4]&p[3]&q[2]  |  p[6]&p[5]&p[4]&p[3]&p[2]&q[1]  |  p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&q[0]  |  p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c0;
         c8  =q[7]  |  p[7]&q[6]  |  p[7]&p[6]&q[5]  |  p[7]&p[6]&p[5]&q[4]  |  p[7]&p[6]&p[5]&p[4]&q[3]  |  p[7]&p[6]&p[5]&p[4]&p[3]&q[2]  |  p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&q[1]  |  p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&q[0]  |  p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&c0;


s[0]=p[0]^q[0]^c0;
s[1]=p[1]^q[1]^c[1];
s[2]=p[2]^q[2]^c[2];
s[3]=p[3]^q[3]^c[3];
s[4]=p[4]^q[4]^c[4];
s[5]=p[5]^q[5]^c[5];
s[6]=p[6]^q[6]^c[6];
s[7]=p[7]^q[7]^c[7];
end

endmodule
