module t_Image_Converter_1(); 
  wire		Done;
  wire 	[1: 8]	HTPV_Row_1, HTPV_Row_2, HTPV_Row_3; 	 
  wire 	[1: 8] 	HTPV_Row_4, HTPV_Row_5, HTPV_Row_6; 

  reg 	[7: 0]	pixel_1,    pixel_2,  pixel_3,   pixel_4,   pixel_5,   pixel_6,   pixel_7,   pixel_8;
  reg	[7: 0]	pixel_9,   pixel_10, pixel_11, pixel_12, pixel_13, pixel_14, pixel_15, pixel_16;
  reg	[7: 0]	pixel_17, pixel_18, pixel_19, pixel_20, pixel_21, pixel_22, pixel_23, pixel_24;
  reg	[7: 0]	pixel_25, pixel_26, pixel_27, pixel_28, pixel_29, pixel_30, pixel_31, pixel_32;
  reg	[7: 0]	pixel_33, pixel_34, pixel_35, pixel_36, pixel_37, pixel_38, pixel_39, pixel_40;
  reg	[7: 0]	pixel_41, pixel_42, pixel_43, pixel_44, pixel_45, pixel_46, pixel_47, pixel_48;
  reg	Go, clk, reset;

Image_Converter_1 M0 ( 
  HTPV_Row_1, HTPV_Row_2, HTPV_Row_3, 	 
  HTPV_Row_4, HTPV_Row_5, HTPV_Row_6, 
  Done,
  pixel_1,    pixel_2,  pixel_3,   pixel_4,   pixel_5,   pixel_6,   pixel_7,   pixel_8,
  pixel_9,   pixel_10, pixel_11, pixel_12, pixel_13, pixel_14, pixel_15, pixel_16,
  pixel_17, pixel_18, pixel_19, pixel_20, pixel_21, pixel_22, pixel_23, pixel_24,
  pixel_25, pixel_26, pixel_27, pixel_28, pixel_29, pixel_30, pixel_31, pixel_32,
  pixel_33, pixel_34, pixel_35, pixel_36, pixel_37, pixel_38, pixel_39, pixel_40,
  pixel_41, pixel_42, pixel_43, pixel_44, pixel_45, pixel_46, pixel_47, pixel_48,
  Go, clk, reset);

initial begin: Image_Pattern_1
    pixel_1 =255;pixel_2 =255;pixel_3 =255;pixel_4 =255;pixel_5 =0;pixel_6 =0;pixel_7 =0;pixel_8 =0;    
    pixel_9 =255; pixel_10 =255; pixel_11 =255;pixel_12 =255;pixel_13 =0;pixel_14 =0;pixel_15 =0;pixel_16 =0;
    pixel_17 =255;pixel_18 =255;pixel_19 =255;pixel_20 =255;pixel_21 =0;pixel_22 =0;pixel_23 =0;pixel_24 =0;
    pixel_25 =0;pixel_26 =0;pixel_27 =0;pixel_28 =0;pixel_29 =255;pixel_30 =255;pixel_31 =255;pixel_32 =255;
    pixel_33 =0;pixel_34 =0;pixel_35 =0;pixel_36 =0;pixel_37 =255;pixel_38 =255;pixel_39 =255;pixel_40 =255;
    pixel_41 =0;pixel_42 =0;pixel_43 =0;pixel_44 =0;pixel_45 =255;pixel_46 =255;pixel_47 =255;pixel_48 =255;
   end

  initial begin: Image_Pattern_2
    #260 
    pixel_1 =0;pixel_2 =0;pixel_3 =0;pixel_4 =0;pixel_5 =255;pixel_6 =255;pixel_7 =255;pixel_8 =255;
    pixel_9 =0;pixel_10 =0;pixel_11 =0;pixel_12 =0;pixel_13 =255;pixel_14 =255;pixel_15 =255;pixel_16 =255;
    pixel_17 =0;pixel_18 =0;pixel_19 =0;pixel_20 =0;pixel_21 =255;pixel_22 =255;pixel_23 =255;pixel_24 =255;
    pixel_25 =255;pixel_26 =255;pixel_27 =255;pixel_28 =255;pixel_29 =0;pixel_30 =0;pixel_31 =0;pixel_32 =0;
    pixel_33 =255;pixel_34 =255;pixel_35 =255;pixel_36 =255;pixel_37 =0;pixel_38 =0;pixel_39 =0;pixel_40 =0;
    pixel_41 =255;pixel_42 =255;pixel_43 =255;pixel_44 =255;pixel_45 =0;pixel_46 =0;pixel_47 =0;pixel_48 =0;
   end

 initial begin: Image_Pattern_3_Cross
    #520
   pixel_1 =0;pixel_2 =0;pixel_3 =255;pixel_4 =255;pixel_5 =255;pixel_6 =255;pixel_7 =0;pixel_8 =0;    
    pixel_9 =0; pixel_10 =0; pixel_11 =255;pixel_12 =255;pixel_13 =255;pixel_14 =255;pixel_15 =0;pixel_16 =0;
    pixel_17 =255;pixel_18 =255;pixel_19 =255;pixel_20 =255;pixel_21 =255;pixel_22 =255;pixel_23 =255;pixel_24 =255;
    pixel_25 =255;pixel_26 =255;pixel_27 =255;pixel_28 =255;pixel_29 =255;pixel_30 =255;pixel_31 =255;pixel_32 =255;
    pixel_33 =0;pixel_34 =0;pixel_35 =255;pixel_36 =255;pixel_37 =255;pixel_38 =255;pixel_39 =0;pixel_40 =0;
    pixel_41 =0;pixel_42 =0;pixel_43 =255;pixel_44 =255;pixel_45 =255;pixel_46 =255;pixel_47 =0;pixel_48 =0;
  end

initial begin: Image_Pattern_4_Bar_Cross  
#780
   pixel_1 =255;pixel_2 =255;pixel_3 =0;pixel_4 =0;pixel_5 =0;pixel_6 =0;pixel_7 =255;pixel_8 =255;    
    pixel_9 =255; pixel_10 =255; pixel_11 =0;pixel_12 =0;pixel_13 =0;pixel_14 =0;pixel_15 =255;pixel_16 =255;
    pixel_17 =255;pixel_18 =255;pixel_19 =255;pixel_20 =255;pixel_21 =255;pixel_22 =255;pixel_23 =255;pixel_24 =255;
    pixel_25 =255;pixel_26 =255;pixel_27 =255;pixel_28 =255;pixel_29 =255;pixel_30 =255;pixel_31 =255;pixel_32 =255;
    pixel_33 =255;pixel_34 =255;pixel_35 =0;pixel_36 =0;pixel_37 =0;pixel_38 =0;pixel_39 =255;pixel_40 =255;
    pixel_41 =255;pixel_42 =255;pixel_43 =0;pixel_44 =0;pixel_45 =0;pixel_46 =0;pixel_47 =255;pixel_48 =255;
  end

  initial begin: Image_Pattern_5_Graduated_Left_to_Right
    #1040    pixel_1 =31;pixel_2 =63;pixel_3 =95;pixel_4 =127;pixel_5 =159;pixel_6 =191;pixel_7 =223;pixel_8 =255;
    pixel_9 =31;pixel_10 =63;pixel_11 =95;pixel_12 =127;pixel_13 =159;pixel_14 =191;pixel_15 =223;pixel_16 =255;
    pixel_17 =31;pixel_18 =63;pixel_19 =95;pixel_20 =127;pixel_21 =159;pixel_22 =191;pixel_23 =223;pixel_24 =255;
    pixel_25 =31;pixel_26 =63;pixel_27 =95;pixel_28 =127;pixel_29 =159;pixel_30 =191;pixel_31 =223;pixel_32 =255;
    pixel_33 =31;pixel_34 =63;pixel_35 =95;pixel_36 =127;pixel_37 =159;pixel_38 =191;pixel_39 =223;pixel_40 =255;
    pixel_41 =31;pixel_42 =63;pixel_43 =95;pixel_44 =127;pixel_45 =159;pixel_46 =191;pixel_47 =223;pixel_48 =255;
  end
  
initial #3200 $finish;
initial begin clk =0; forever #5 clk = ~clk; end

  initial fork
    #10 reset= 1; 
    #30 reset = 0; 
  join

  initial fork
    #50 Go = 1; 		// Image #1
    #60 Go = 0;
 
    #270 reset = 1;		// Image #2
    #290 reset = 0;
   #300 Go = 1;
   #310 Go = 0;

    #600 reset = 1;		// Image #3
    #630 reset = 0;
    #680 Go = 1;
    #690 Go = 0;

    #900 reset = 1;		// Image #4
    #930 reset = 0;
    #980 Go = 1;
    #990 Go = 0;

    #1200 reset = 1;	// Image #5
    #1230 reset = 0;
    #1280 Go = 1;
    #1290 Go = 0;
  join
endmodule

